version https://git-lfs.github.com/spec/v1
oid sha256:7ef49a47c227ccdee67a19c33777fe3308251eb53dc87a172662d42690741a8a
size 17951748
