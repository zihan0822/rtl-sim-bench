version https://git-lfs.github.com/spec/v1
oid sha256:e726455d8cd87cacf1f0d3037cdb6758b1282c1766ad50ef57428a3ae7036c5a
size 4119656
