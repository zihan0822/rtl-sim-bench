version https://git-lfs.github.com/spec/v1
oid sha256:0aa0f78f2e9fbf74d16c3e5aaa1aba0329681bb7599bf79a3a514239dc43ba90
size 17951237
