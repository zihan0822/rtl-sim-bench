version https://git-lfs.github.com/spec/v1
oid sha256:8f103a7d94dcacea71fa84e9e1b6e8471c91efdc513f038d242c13de5420297e
size 4118388
